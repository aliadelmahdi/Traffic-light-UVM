module golden_model(
 
);

  

endmodule