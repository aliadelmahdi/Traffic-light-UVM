`include "traffic_light_defines.svh" // For macros
`timescale `TIME_UNIT / `TIME_PRECISION

module traffic_light_sva(

  );
 
endmodule


