interface traffic_if(input bit clk);
   
endinterface
